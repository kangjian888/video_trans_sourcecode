`timescales 1ns/1ps

module(
	);
reg clk, reset, 
    
endmodule